library ieee;
context ieee.ieee_std_context;
use ieee.math_real.all;

library std;
use std.textio.all;

entity testbench is
end entity testbench;

architecture rtl of testbench is

begin

	

end architecture;