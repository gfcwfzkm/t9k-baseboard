library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity top is
	port (
		clk   : in std_logic;
		reset : in std_logic		
	);
end entity top;

architecture rtl of top is

begin

	

end architecture;